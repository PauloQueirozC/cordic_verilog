module negacao(input [3:0] A, output [3:0] B);
	assign B = -A;
endmodule